`timescale 10ns/10ps
module full_tb;
reg a,b,cin;
wire sum,cout;
full_adder ga(a,b,cin,sum,cout);
initial begin
a=0;b=0;cin=0;
#10 a=0;b=1;cin=0;
#10 a=0;b=0;cin=1;
#10 a=1;b=0;cin=0;
#10 a=1;b=0;cin=1;
#10 a=1;b=1;cin=0;
#10 a=1;b=1;cin=1;
#40;
end
endmodule

